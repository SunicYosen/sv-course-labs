`ifndef INC_SCOREBOARD_SV
`define INC_SCOREBOARD_SV
class Scoreboard;
//  extern function new(string name = "Scoreboard", pkt_mbox driver_mbox = null, receiver_mbox = null);
//  extern virtual function void check();           //Compare the data package and check the correctness
endclass: Scoreboard

`endif

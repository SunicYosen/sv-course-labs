`ifndef INC_RECEIVERBASE_SV
`define INC_RECEIVERBASE_SV
class Receiver;
//   extern function new(string name = "ReceiverBase", virtual router_io.TB rtr_io);
//   extern virtual  task recv();    // Receive packets from the DUT output port
endclass
`endif
